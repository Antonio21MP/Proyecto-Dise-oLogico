`timescale 1ns / 1ps
module LEDS_CONTROL(
	input 
	output
    );


endmodule
